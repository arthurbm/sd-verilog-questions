module mux4_to_1 (
    output wire F,
    input wire A, B, C, D, E, F
);
    
endmodule